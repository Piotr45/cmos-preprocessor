.subckt DIODA in vss vdd
Mn0 in in VSS VSS nch w=0.3u l=0.44u
Mp0 in in VDD VDD pch w=1.715u l=0.44u
.ends DIODA
