*** PREPROCESSOR
.INCLUDE components/AXON.sp
.INCLUDE components/DENDRITE.sp
.INCLUDE components/CMRR.sp

.subckt PREPROCESSOR IN0p IN0m IN1p IN1m OUT0p OUT0m VSS VDD

xCMp_0 IN0p OUTn_n1p0 OUTn_n2p0 VSS VDD CM2
xCMm_0 IN0m OUTp_n1p0 OUTp_n2p0 VSS VDD CM2
xCMp_1 IN1p OUTn_n1p1 OUTn_n2p1 VSS VDD CM2
xCMm_1 IN1m OUTp_n1p1 OUTp_n2p1 VSS VDD CM2

xDENDRYTw0n0d0 OUTn_n1p0 OUTp_n1p0 OUTmw0_n0 OUTpw0_n0 VDD VSS VDD VDD VDD VSS VDD VSS VSS VSS VSS VSS VSS VDD DENDRYT
xDENDRYTw0n0d1 OUTp_n1p0 OUTn_n1p0 OUTmw0_n0 OUTpw0_n0 VSS VSS VSS VSS VDD VSS VDD VDD VDD VDD VDD VDD VSS VDD DENDRYT

xDENDRYTw0n1d0 OUTn_n1p1 OUTp_n1p1 OUTmw0_n1 OUTpw0_n1 VDD VSS VDD VDD VDD VSS VDD VSS VDD VSS VDD VDD VSS VDD DENDRYT
xDENDRYTw0n1d1 OUTn_n1p1 OUTp_n1p1 OUTmw0_n1 OUTpw0_n1 VSS VDD VSS VDD VDD VSS VDD VDD VDD VSS VSS VSS VSS VDD DENDRYT

xAKSONw0n0 OUTpw0_n0 OUTmw0_n0 OUTp_w0n0 OUTm_w0n0 VSS VDD AKSON
xAKSONw0n1 OUTpw0_n1 OUTmw0_n1 OUTp_w0n1 OUTm_w0n1 VSS VDD AKSON

xCMRRw0n0 OUTp_w0n0 OUTm_w0n0 INw2p_n1p0 INw2m_n1p0 VSS VDD CMRR
xCMRRw0n1 OUTp_w0n1 OUTm_w0n1 INw2p_n1p1 INw2m_n1p1 VSS VDD CMRR

xDENDRYTw1n0d0 OUTn_n1p0 OUTp_n1p0 OUTmw1_n0 OUTpw1_n0 VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VSS VDD VSS VDD DENDRYT

xAKSONw1n0 OUTpw1_n0 OUTmw1_n0 OUTp_w1n0 OUTm_w1n0 VSS VDD AKSON

xCMRRw1n0 OUTp_w1n0 OUTm_w1n0 OUT0p OUT0m VSS VDD CMRR

.ends PREPROCESSOR